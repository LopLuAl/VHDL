LED 0 50 Hz TODOS LOS DUTY
01000001 00000000   
01000001 00000001 
01000001 00000010 
01000001 00000011
LED 1 80 Hz TODOS LOS DUTY
01000001 01010000
01000001 01010001
01000001 01010010
01000001 01010011
LED 2 100 Hz TODOS LOS DUTY
01000001 10100000
01000001 10100001
01000001 10100010
01000001 10100011
LED 3 125 Hz TODOS LOS DUTY
01000001 11110000
01000001 11110001
01000001 11110010
01000001 11110011